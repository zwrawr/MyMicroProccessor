
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity register is
    Port ( clk : in  STD_LOGIC;
           data_in : in  STD_LOGIC_VECTOR (3 downto 0);
           data_out : out  STD_LOGIC_VECTOR (3 downto 0));
end register;

architecture Behavioral of register is

begin


end Behavioral;

